    Mac OS X            	   2         �                                      ATTR       �   �                     �     com.dropbox.attrs    

��i��N<     |`h莄