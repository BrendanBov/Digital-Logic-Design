module control();
//State machine in top.sv
endmodule
